class simple_sequencer extends uvm_sequencer #(simple_item, simple_rsp);


endclass
